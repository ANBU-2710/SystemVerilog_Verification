class transaction;
  
  rand bit a,b,c_in;
  bit sum,c_out;
  
endclass